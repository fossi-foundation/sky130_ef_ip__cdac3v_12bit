magic
tech sky130A
magscale 1 2
timestamp 1747669346
<< nwell >>
rect 58549 -26640 83864 21013
<< mvnsubdiff >>
rect 58615 20927 83798 20947
rect 58615 20893 58695 20927
rect 83718 20893 83798 20927
rect 58615 20873 83798 20893
rect 58615 20867 58689 20873
rect 58615 -26494 58635 20867
rect 58669 -26494 58689 20867
rect 58615 -26500 58689 -26494
rect 83724 20867 83798 20873
rect 83724 -26494 83744 20867
rect 83778 -26494 83798 20867
rect 83724 -26500 83798 -26494
rect 58615 -26520 83798 -26500
rect 58615 -26554 58695 -26520
rect 83718 -26554 83798 -26520
rect 58615 -26574 83798 -26554
<< mvnsubdiffcont >>
rect 58695 20893 83718 20927
rect 58635 -26494 58669 20867
rect 83744 -26494 83778 20867
rect 58695 -26554 83718 -26520
<< locali >>
rect 58615 20927 83798 20947
rect 58615 20893 58695 20927
rect 83718 20893 83798 20927
rect 58615 20873 83798 20893
rect 58615 20867 58689 20873
rect 58615 -26494 58635 20867
rect 58669 -26494 58689 20867
rect 58615 -26500 58689 -26494
rect 83724 20867 83798 20873
rect 83724 -26494 83744 20867
rect 83778 -26494 83798 20867
rect 83724 -26500 83798 -26494
rect 58615 -26520 83798 -26500
rect 58615 -26554 58695 -26520
rect 83718 -26554 83798 -26520
rect 58615 -26574 83798 -26554
<< metal3 >>
rect 58361 18300 58817 18364
rect 83378 18176 83379 18240
rect 83445 18176 83446 18240
rect 83523 18176 84124 18240
rect 58323 15820 58917 15884
rect 58987 15820 58988 15884
rect 59052 15820 59053 15884
rect 83503 15696 83504 15760
rect 83568 15696 83569 15760
rect 58865 13340 58866 13404
rect 58930 13340 58931 13404
rect 83378 13216 83379 13280
rect 83445 13216 83446 13280
rect 58988 10860 58989 10924
rect 59053 10860 59054 10924
rect 58342 10736 58743 10800
rect 58807 10736 58980 10800
rect 81945 10546 82005 10770
rect 58865 8380 58866 8444
rect 58930 8380 58931 8444
rect 83445 8256 83997 8320
rect 58737 5900 58743 5964
rect 58807 5900 58879 5964
rect 58988 5776 58989 5840
rect 59053 5776 59054 5840
rect 83378 3420 83379 3484
rect 83445 3420 83446 3484
rect 58256 3296 58866 3360
rect 58930 3296 59007 3360
rect 83448 940 83504 1004
rect 83568 940 83982 1004
rect 83534 -1664 84044 -1600
rect 69804 -4031 69860 -3967
rect 70081 -4031 70102 -3967
rect 83551 -4031 84044 -3967
rect 58988 -4155 58989 -4091
rect 59053 -4155 59054 -4091
rect 83379 -6511 83380 -6447
rect 83444 -6511 83445 -6447
rect 58306 -6635 58866 -6571
rect 58930 -6635 58989 -6571
rect 83454 -8991 83503 -8927
rect 83567 -8991 84023 -8927
rect 58988 -9115 58989 -9051
rect 59053 -9115 59054 -9051
rect 83379 -11471 83380 -11407
rect 83444 -11471 83445 -11407
rect 83551 -11595 83626 -11531
rect 83690 -11595 83700 -11531
rect 58383 -13951 58879 -13887
rect 83502 -14075 83503 -14011
rect 83567 -14075 83568 -14011
rect 58346 -16431 58879 -16367
rect 83551 -16431 83626 -16367
rect 83690 -16431 84056 -16367
rect 83379 -16555 83380 -16491
rect 83444 -16555 83445 -16491
rect 58988 -18911 58989 -18847
rect 59053 -18911 59054 -18847
rect 58865 -21391 58866 -21327
rect 58930 -21391 58931 -21327
rect 83379 -21515 83380 -21451
rect 83444 -21515 83445 -21451
rect 83514 -21515 84033 -21451
rect 58243 -23871 58911 -23807
rect 83610 -23995 84044 -23931
<< via3 >>
rect 83379 18176 83445 18240
rect 58988 15820 59052 15884
rect 83504 15696 83568 15760
rect 58866 13340 58930 13404
rect 83379 13216 83445 13280
rect 58989 10860 59053 10924
rect 58743 10736 58807 10800
rect 72347 10736 72565 10800
rect 58866 8380 58930 8444
rect 58743 5900 58807 5964
rect 58989 5776 59053 5840
rect 83379 3420 83445 3484
rect 58866 3296 58930 3360
rect 83504 940 83568 1004
rect 58989 816 59053 880
rect 83379 -1540 83445 -1476
rect 69860 -1664 70081 -1600
rect 69860 -4031 70081 -3967
rect 58989 -4155 59053 -4091
rect 83380 -6511 83444 -6447
rect 58866 -6635 58930 -6571
rect 83503 -8991 83567 -8927
rect 58989 -9115 59053 -9051
rect 83380 -11471 83444 -11407
rect 83626 -11595 83690 -11531
rect 83503 -14075 83567 -14011
rect 83626 -16431 83690 -16367
rect 83380 -16555 83444 -16491
rect 58989 -18911 59053 -18847
rect 83503 -19035 83567 -18971
rect 58866 -21391 58930 -21327
rect 83380 -21515 83444 -21451
rect 58989 -23871 59053 -23807
<< metal4 >>
rect 83382 18241 83442 18381
rect 83378 18240 83446 18241
rect 83378 18176 83379 18240
rect 83445 18176 83446 18240
rect 83378 18175 83446 18176
rect 58991 15885 59051 15918
rect 58987 15884 59053 15885
rect 58987 15820 58988 15884
rect 59052 15820 59053 15884
rect 58987 15819 59053 15820
rect 58868 13405 58928 13452
rect 58865 13404 58931 13405
rect 58865 13340 58866 13404
rect 58930 13340 58931 13404
rect 58865 13339 58931 13340
rect 58745 10801 58805 10812
rect 58742 10800 58808 10801
rect 58742 10736 58743 10800
rect 58807 10736 58808 10800
rect 58742 10735 58808 10736
rect 58745 5965 58805 10735
rect 58868 8445 58928 13339
rect 58991 10925 59051 15819
rect 83382 13281 83442 18175
rect 83506 15761 83566 15781
rect 83503 15760 83569 15761
rect 83503 15696 83504 15760
rect 83568 15696 83569 15760
rect 83503 15695 83569 15696
rect 83378 13280 83446 13281
rect 83378 13216 83379 13280
rect 83445 13216 83446 13280
rect 83378 13215 83446 13216
rect 58988 10924 59054 10925
rect 58988 10860 58989 10924
rect 59053 10860 59054 10924
rect 58988 10859 59054 10860
rect 58865 8444 58931 8445
rect 58865 8380 58866 8444
rect 58930 8380 58931 8444
rect 58865 8379 58931 8380
rect 58742 5964 58808 5965
rect 58742 5900 58743 5964
rect 58807 5900 58808 5964
rect 58742 5899 58808 5900
rect 58745 5867 58805 5899
rect 58868 3361 58928 8379
rect 58991 5841 59051 10859
rect 72346 10800 72566 10801
rect 72346 10736 72347 10800
rect 72565 10736 72566 10800
rect 72346 10735 72566 10736
rect 72425 10470 72485 10735
rect 58988 5840 59054 5841
rect 58988 5776 58989 5840
rect 59053 5776 59054 5840
rect 58988 5775 59054 5776
rect 58865 3360 58931 3361
rect 58865 3296 58866 3360
rect 58930 3296 58931 3360
rect 58865 3295 58931 3296
rect 58868 3268 58928 3295
rect 58991 881 59051 5775
rect 83382 3485 83442 13215
rect 83378 3484 83446 3485
rect 83378 3420 83379 3484
rect 83445 3420 83446 3484
rect 83378 3419 83446 3420
rect 58988 880 59054 881
rect 58988 816 58989 880
rect 59053 816 59054 880
rect 58988 815 59054 816
rect 58991 786 59051 815
rect 60025 -1930 60085 -1210
rect 69945 -1599 70005 -1150
rect 69859 -1600 70082 -1599
rect 69859 -1664 69860 -1600
rect 70081 -1664 70082 -1600
rect 69859 -1665 70082 -1664
rect 82345 -1930 82405 -1210
rect 83382 -1475 83442 3419
rect 83506 1005 83566 15695
rect 83503 1004 83569 1005
rect 83503 940 83504 1004
rect 83568 940 83569 1004
rect 83503 939 83569 940
rect 83506 929 83566 939
rect 83378 -1476 83446 -1475
rect 83378 -1540 83379 -1476
rect 83445 -1540 83446 -1476
rect 83378 -1541 83446 -1540
rect 83382 -1564 83442 -1541
rect 60935 -2845 61655 -2785
rect 63415 -2845 64135 -2785
rect 65895 -2845 66615 -2785
rect 73335 -2845 74055 -2785
rect 75815 -2845 76535 -2785
rect 78295 -2845 79015 -2785
rect 80775 -2845 81495 -2785
rect 58991 -4090 59051 -4066
rect 58988 -4091 59054 -4090
rect 58988 -4155 58989 -4091
rect 59053 -4155 59054 -4091
rect 58988 -4156 59054 -4155
rect 58868 -6570 58928 -6535
rect 58865 -6571 58931 -6570
rect 58865 -6635 58866 -6571
rect 58930 -6635 58931 -6571
rect 58865 -6636 58931 -6635
rect 58868 -21326 58928 -6636
rect 58991 -9050 59051 -4156
rect 60025 -4421 60085 -3701
rect 69945 -3966 70005 -3700
rect 69859 -3967 70082 -3966
rect 69859 -4031 69860 -3967
rect 70081 -4031 70082 -3967
rect 69859 -4032 70082 -4031
rect 69945 -4421 70005 -4032
rect 82345 -4421 82405 -3701
rect 83382 -6446 83442 -6397
rect 83379 -6447 83445 -6446
rect 83379 -6511 83380 -6447
rect 83444 -6511 83445 -6447
rect 83379 -6512 83445 -6511
rect 58988 -9051 59054 -9050
rect 58988 -9115 58989 -9051
rect 59053 -9115 59054 -9051
rect 58988 -9116 59054 -9115
rect 58991 -18846 59051 -9116
rect 83382 -11406 83442 -6512
rect 83505 -8926 83565 -8915
rect 83502 -8927 83568 -8926
rect 83502 -8991 83503 -8927
rect 83567 -8991 83568 -8927
rect 83502 -8992 83568 -8991
rect 83379 -11407 83445 -11406
rect 83379 -11471 83380 -11407
rect 83444 -11471 83445 -11407
rect 83379 -11472 83445 -11471
rect 69945 -14341 70005 -13621
rect 68375 -15251 69095 -15191
rect 70855 -15251 71575 -15191
rect 69945 -16821 70005 -16101
rect 83382 -16490 83442 -11472
rect 83505 -14010 83565 -8992
rect 83628 -11530 83688 -11496
rect 83625 -11531 83691 -11530
rect 83625 -11595 83626 -11531
rect 83690 -11595 83691 -11531
rect 83625 -11596 83691 -11595
rect 83502 -14011 83568 -14010
rect 83502 -14075 83503 -14011
rect 83567 -14075 83568 -14011
rect 83502 -14076 83568 -14075
rect 83379 -16491 83445 -16490
rect 83379 -16555 83380 -16491
rect 83444 -16555 83445 -16491
rect 83379 -16556 83445 -16555
rect 58988 -18847 59054 -18846
rect 58988 -18911 58989 -18847
rect 59053 -18911 59054 -18847
rect 58988 -18912 59054 -18911
rect 58865 -21327 58931 -21326
rect 58865 -21391 58866 -21327
rect 58930 -21391 58931 -21327
rect 58865 -21392 58931 -21391
rect 58868 -21562 58928 -21392
rect 58991 -23806 59051 -18912
rect 83382 -21450 83442 -16556
rect 83505 -18970 83565 -14076
rect 83628 -16366 83688 -11596
rect 83625 -16367 83691 -16366
rect 83625 -16431 83626 -16367
rect 83690 -16431 83691 -16367
rect 83625 -16432 83691 -16431
rect 83628 -16450 83688 -16432
rect 83502 -18971 83568 -18970
rect 83502 -19035 83503 -18971
rect 83567 -19035 83568 -18971
rect 83502 -19036 83568 -19035
rect 83505 -19061 83565 -19036
rect 83379 -21451 83445 -21450
rect 83379 -21515 83380 -21451
rect 83444 -21515 83445 -21451
rect 83379 -21516 83445 -21515
rect 83382 -21534 83442 -21516
rect 58988 -23807 59054 -23806
rect 58988 -23871 58989 -23807
rect 59053 -23871 59054 -23807
rect 58988 -23872 59054 -23871
rect 58991 -24038 59051 -23872
use cap_array_half  cap_array_half_0
timestamp 1747669346
transform -1 0 164043 0 -1 -5787
box 80293 -26673 105363 -4081
use cap_array_half  cap_array_half_1
timestamp 1747669346
transform 1 0 -21613 0 1 156
box 80293 -26673 105363 -4081
use caparray_connect_near  caparray_connect_near_0
timestamp 1747669346
transform -1 0 151643 0 -1 -28107
box 80427 -26673 82908 -26177
use cdac_cross2_short  cdac_cross2_short_0
timestamp 1747669346
transform 1 0 14880 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_1
timestamp 1747669346
transform 1 0 -4960 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_2
timestamp 1747669346
transform 1 0 -2480 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_3
timestamp 1747669346
transform 1 0 0 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_6
timestamp 1747669346
transform 1 0 7440 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_7
timestamp 1747669346
transform 1 0 9920 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross2_short  cdac_cross2_short_8
timestamp 1747669346
transform 1 0 12400 0 1 0
box 65895 -3386 66615 -2244
use cdac_cross_short  cdac_cross_short_0
timestamp 1747669346
transform 0 1 62881 -1 0 64685
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_1
timestamp 1747669346
transform 1 0 14880 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_2
timestamp 1747669346
transform 1 0 -4960 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_3
timestamp 1747669346
transform 1 0 -2480 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_4
timestamp 1747669346
transform 1 0 0 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_5
timestamp 1747669346
transform 1 0 2480 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_6
timestamp 1747669346
transform 1 0 4960 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_7
timestamp 1747669346
transform 1 0 7440 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_8
timestamp 1747669346
transform 1 0 9920 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_9
timestamp 1747669346
transform 1 0 12400 0 1 -22315
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_10
timestamp 1747669346
transform 0 -1 57229 1 0 -75276
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_11
timestamp 1747669346
transform 0 -1 57229 1 0 -77756
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_12
timestamp 1747669346
transform 0 -1 57229 1 0 -87676
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_13
timestamp 1747669346
transform 0 -1 57229 1 0 -82716
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_14
timestamp 1747669346
transform 0 -1 57229 1 0 -85196
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_15
timestamp 1747669346
transform 0 1 62881 -1 0 82045
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_16
timestamp 1747669346
transform 0 1 85201 -1 0 82045
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_17
timestamp 1747669346
transform 0 1 85201 -1 0 47314
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_18
timestamp 1747669346
transform 0 1 85201 -1 0 49794
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_19
timestamp 1747669346
transform 0 1 85201 -1 0 52274
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_20
timestamp 1747669346
transform 0 1 85201 -1 0 54754
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_21
timestamp 1747669346
transform 0 1 85201 -1 0 57234
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_22
timestamp 1747669346
transform 0 1 85201 -1 0 59714
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_23
timestamp 1747669346
transform 0 1 85201 -1 0 62194
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_24
timestamp 1747669346
transform 0 1 85201 -1 0 64685
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_25
timestamp 1747669346
transform 0 1 85201 -1 0 67165
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_26
timestamp 1747669346
transform 0 1 85201 -1 0 69645
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_27
timestamp 1747669346
transform 0 1 85201 -1 0 72125
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_28
timestamp 1747669346
transform 0 1 85201 -1 0 74605
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_29
timestamp 1747669346
transform 0 1 85201 -1 0 77085
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_30
timestamp 1747669346
transform 0 1 85201 -1 0 79565
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_31
timestamp 1747669346
transform 0 1 85201 -1 0 44834
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_32
timestamp 1747669346
transform 0 -1 57229 1 0 -80236
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_33
timestamp 1747669346
transform 0 -1 57229 1 0 -72796
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_34
timestamp 1747669346
transform 0 -1 57229 1 0 -70316
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_35
timestamp 1747669346
transform 0 1 62881 -1 0 72125
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_36
timestamp 1747669346
transform 0 1 62881 -1 0 69645
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_37
timestamp 1747669346
transform 0 1 62881 -1 0 67165
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_38
timestamp 1747669346
transform 0 1 62881 -1 0 79565
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_39
timestamp 1747669346
transform 0 1 62881 -1 0 77085
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_40
timestamp 1747669346
transform 0 1 62881 -1 0 74605
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_41
timestamp 1747669346
transform 1 0 14880 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_42
timestamp 1747669346
transform 1 0 12400 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_43
timestamp 1747669346
transform 1 0 9920 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_44
timestamp 1747669346
transform 1 0 7440 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_45
timestamp 1747669346
transform 1 0 4960 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_46
timestamp 1747669346
transform 1 0 2480 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_47
timestamp 1747669346
transform 1 0 0 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_48
timestamp 1747669346
transform 1 0 -2480 0 1 22336
box 65895 -3386 66615 -2266
use cdac_cross_short  cdac_cross_short_49
timestamp 1747669346
transform 1 0 -4960 0 1 22336
box 65895 -3386 66615 -2266
use cdac_ratioed_cap  cdac_ratioed_cap_0
array 0 9 2480 0 0 2797
timestamp 1747669346
transform 1 0 -21716 0 1 29649
box 80396 -33846 83146 -31084
<< labels >>
flabel comment 58859 -4132 58859 -4132 0 FreeSans 800 0 0 0 D4
flabel comment 83585 -1497 83585 -1497 0 FreeSans 800 0 0 0 D10
flabel metal3 58308 -6635 58508 -6571 0 FreeSans 480 0 0 0 D2
port 8 nsew
flabel metal3 58386 -13951 58545 -13887 0 FreeSans 480 0 0 0 D0
port 1 nsew
flabel metal3 58244 -23871 58444 -23807 0 FreeSans 480 0 0 0 D4
port 2 nsew
flabel metal3 83830 -21515 84030 -21451 0 FreeSans 480 0 0 0 D5
port 5 nsew
flabel metal3 83854 -16431 84054 -16367 0 FreeSans 480 0 0 0 D1
port 6 nsew
flabel metal3 83822 -8991 84022 -8927 0 FreeSans 480 0 0 0 D3
port 12 nsew
flabel metal4 83544 -16396 83544 -16396 0 FreeSans 800 0 0 0 D1
flabel comment 83563 -6484 83563 -6484 0 FreeSans 800 0 0 0 D5
flabel metal4 83563 -11436 83563 -11436 0 FreeSans 800 0 0 0 D5
flabel metal4 83563 -16519 83563 -16519 0 FreeSans 800 0 0 0 D5
flabel metal3 83574 -21477 83574 -21477 0 FreeSans 800 0 0 0 D5
flabel metal3 83579 -8963 83579 -8963 0 FreeSans 800 0 0 0 D3
flabel comment 83584 -14047 83584 -14047 0 FreeSans 800 0 0 0 D3
flabel comment 83582 -19005 83582 -19005 0 FreeSans 800 0 0 0 D3
flabel metal3 83576 -11564 83576 -11564 0 FreeSans 800 0 0 0 D1
flabel metal4 58868 -11565 58868 -11565 0 FreeSans 800 0 0 0 D1
flabel metal4 58877 -13917 58877 -13917 0 FreeSans 800 0 0 0 D0
flabel comment 58859 -9078 58859 -9078 0 FreeSans 800 0 0 0 D4
flabel comment 58864 -18878 58864 -18878 0 FreeSans 800 0 0 0 D4
flabel metal3 58850 -23844 58850 -23844 0 FreeSans 800 0 0 0 D4
flabel metal3 58858 -6605 58858 -6605 0 FreeSans 800 0 0 0 D2
flabel comment 58853 -21361 58853 -21361 0 FreeSans 800 0 0 0 D2
flabel metal3 83840 -4031 84040 -3967 0 FreeSans 480 0 0 0 VP1
port 3 nsew
flabel metal3 58344 10736 58544 10800 0 FreeSans 480 0 0 0 D7
port 11 nsew
flabel metal3 58258 3296 58458 3360 0 FreeSans 480 0 0 0 D9
port 4 nsew
flabel metal3 58324 15820 58516 15884 0 FreeSans 480 0 0 0 D11
port 14 nsew
flabel metal3 83780 940 83980 1004 0 FreeSans 480 0 0 0 D8
port 0 nsew
flabel metal3 83798 8256 83997 8320 0 FreeSans 480 0 0 0 D6
port 9 nsew
flabel metal3 83928 18176 84120 18240 0 FreeSans 480 0 0 0 D10
port 13 nsew
flabel metal4 83561 3454 83561 3454 0 FreeSans 800 0 0 0 D10
flabel metal3 83572 18206 83572 18206 0 FreeSans 800 0 0 0 D10
flabel comment 83568 13247 83568 13247 0 FreeSans 800 0 0 0 D10
flabel comment 83573 15730 83573 15730 0 FreeSans 800 0 0 0 D8
flabel metal3 83584 971 83584 971 0 FreeSans 800 0 0 0 D8
flabel metal3 83572 8289 83572 8289 0 FreeSans 800 0 0 0 D6
flabel comment 83580 10769 83580 10769 0 FreeSans 800 0 0 0 VSS
flabel metal3 58859 15856 58859 15856 0 FreeSans 800 0 0 0 D11
flabel comment 58855 10886 58855 10886 0 FreeSans 800 0 0 0 D11
flabel comment 58855 5807 58855 5807 0 FreeSans 800 0 0 0 D11
flabel comment 58855 845 58855 845 0 FreeSans 800 0 0 0 D11
flabel comment 58859 13369 58859 13369 0 FreeSans 800 0 0 0 D9
flabel comment 58843 8408 58843 8408 0 FreeSans 800 0 0 0 D9
flabel metal3 58837 3316 58837 3316 0 FreeSans 800 0 0 0 D9
flabel metal3 58847 10760 58847 10760 0 FreeSans 800 0 0 0 D7
flabel metal3 58847 5928 58847 5928 0 FreeSans 800 0 0 0 D7
flabel metal3 83848 -1664 84044 -1600 0 FreeSans 480 0 0 0 VP2
port 7 nsew
flabel metal4 58889 -16197 58889 -16197 0 FreeSans 800 0 0 0 VSS
flabel metal3 83846 -23995 84043 -23931 0 FreeSans 480 0 0 0 VSS
port 10 nsew
flabel metal3 58346 -16431 58512 -16367 0 FreeSans 480 0 0 0 Vref
port 15 nsew
<< end >>
