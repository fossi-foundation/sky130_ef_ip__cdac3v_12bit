magic
tech sky130A
magscale 1 2
timestamp 1747671550
<< dnwell >>
rect 44121 -15586 48345 -14252
<< nwell >>
rect 44011 -14464 48454 -14149
rect 44011 -15380 46465 -14464
rect 48139 -15380 48454 -14464
rect 44011 -15695 48454 -15380
<< pwell >>
rect 46546 -15380 48139 -14464
<< mvpsubdiff >>
rect 46582 -14564 48050 -14552
rect 46582 -14598 46690 -14564
rect 46958 -14598 47106 -14564
rect 47532 -14598 47680 -14564
rect 47948 -14598 48050 -14564
rect 46582 -14610 48050 -14598
rect 46582 -14638 46640 -14610
rect 46582 -15206 46594 -14638
rect 46628 -15206 46640 -14638
rect 46582 -15234 46640 -15206
rect 46998 -14638 47056 -14610
rect 46998 -15206 47010 -14638
rect 47044 -15206 47056 -14638
rect 46998 -15234 47056 -15206
rect 47572 -14638 47630 -14610
rect 47572 -15206 47584 -14638
rect 47618 -15206 47630 -14638
rect 47572 -15234 47630 -15206
rect 47992 -14638 48050 -14610
rect 47992 -15206 48004 -14638
rect 48038 -15206 48050 -14638
rect 47992 -15234 48050 -15206
rect 46582 -15246 48050 -15234
rect 46582 -15280 46690 -15246
rect 46958 -15280 47106 -15246
rect 47532 -15280 47680 -15246
rect 47948 -15280 48050 -15246
rect 46582 -15292 48050 -15280
<< mvnsubdiff >>
rect 44078 -14235 48388 -14215
rect 44078 -14269 44158 -14235
rect 48308 -14269 48388 -14235
rect 44078 -14289 48388 -14269
rect 44078 -14295 44152 -14289
rect 44078 -15549 44098 -14295
rect 44132 -15549 44152 -14295
rect 48314 -14295 48388 -14289
rect 44273 -14514 46399 -14502
rect 44273 -14548 44381 -14514
rect 44807 -14548 44965 -14514
rect 45463 -14548 45803 -14514
rect 46291 -14548 46399 -14514
rect 44273 -14560 46399 -14548
rect 44273 -14610 44331 -14560
rect 44273 -15256 44285 -14610
rect 44319 -15256 44331 -14610
rect 44273 -15306 44331 -15256
rect 44857 -14610 44915 -14560
rect 44857 -15256 44869 -14610
rect 44903 -15256 44915 -14610
rect 44857 -15306 44915 -15256
rect 45757 -14610 45815 -14560
rect 45757 -15256 45769 -14610
rect 45803 -15256 45815 -14610
rect 45757 -15306 45815 -15256
rect 46341 -14610 46399 -14560
rect 46341 -15256 46353 -14610
rect 46387 -15256 46399 -14610
rect 46341 -15306 46399 -15256
rect 44273 -15318 46399 -15306
rect 44273 -15352 44381 -15318
rect 45707 -15352 45865 -15318
rect 46291 -15352 46399 -15318
rect 44273 -15364 46399 -15352
rect 44078 -15555 44152 -15549
rect 48314 -15549 48334 -14295
rect 48368 -15549 48388 -14295
rect 48314 -15555 48388 -15549
rect 44078 -15575 48388 -15555
rect 44078 -15609 44158 -15575
rect 48308 -15609 48388 -15575
rect 44078 -15629 48388 -15609
<< mvpsubdiffcont >>
rect 46690 -14598 46958 -14564
rect 47106 -14598 47532 -14564
rect 47680 -14598 47948 -14564
rect 46594 -15206 46628 -14638
rect 47010 -15206 47044 -14638
rect 47584 -15206 47618 -14638
rect 48004 -15206 48038 -14638
rect 46690 -15280 46958 -15246
rect 47106 -15280 47532 -15246
rect 47680 -15280 47948 -15246
<< mvnsubdiffcont >>
rect 44158 -14269 48308 -14235
rect 44098 -15549 44132 -14295
rect 44381 -14548 44807 -14514
rect 44965 -14548 45463 -14514
rect 45803 -14548 46291 -14514
rect 44285 -15256 44319 -14610
rect 44869 -15256 44903 -14610
rect 45769 -15256 45803 -14610
rect 46353 -15256 46387 -14610
rect 44381 -15352 45707 -15318
rect 45865 -15352 46291 -15318
rect 48334 -15549 48368 -14295
rect 44158 -15609 48308 -15575
<< locali >>
rect 44098 -14269 44158 -14235
rect 48308 -14269 48368 -14235
rect 44098 -14295 48368 -14269
rect 44132 -14369 48334 -14295
rect 44132 -14514 44319 -14369
rect 46594 -14467 48071 -14449
rect 46594 -14504 46637 -14467
rect 47854 -14504 48071 -14467
rect 44132 -14548 44381 -14514
rect 44807 -14548 44965 -14514
rect 45463 -14548 45803 -14514
rect 46291 -14548 46387 -14514
rect 44132 -14610 44319 -14548
rect 44132 -15256 44285 -14610
rect 44132 -15294 44319 -15256
rect 44869 -14610 44903 -14548
rect 44869 -15294 44903 -15256
rect 45769 -14610 45803 -14548
rect 45769 -15294 45803 -15256
rect 46353 -14610 46387 -14548
rect 46353 -15294 46387 -15256
rect 46594 -14564 48071 -14504
rect 46594 -14598 46690 -14564
rect 46958 -14598 47106 -14564
rect 47532 -14598 47680 -14564
rect 47948 -14598 48071 -14564
rect 46594 -14618 48071 -14598
rect 46594 -14638 46628 -14618
rect 46594 -15246 46628 -15206
rect 47010 -14638 47044 -14618
rect 47010 -15246 47044 -15206
rect 47584 -14638 47618 -14618
rect 47584 -15246 47618 -15206
rect 48004 -14638 48038 -14618
rect 48004 -15246 48038 -15206
rect 46594 -15280 46690 -15246
rect 46958 -15280 47106 -15246
rect 47532 -15280 47680 -15246
rect 47948 -15280 48038 -15246
rect 44132 -15318 46388 -15294
rect 44132 -15352 44381 -15318
rect 45707 -15345 45865 -15318
rect 46291 -15345 46388 -15318
rect 44132 -15380 44500 -15352
rect 46363 -15380 46388 -15345
rect 44132 -15388 46388 -15380
rect 46594 -15355 48036 -15280
rect 44132 -15473 44319 -15388
rect 46594 -15401 46616 -15355
rect 48018 -15401 48036 -15355
rect 46594 -15411 48036 -15401
rect 48210 -15473 48334 -14369
rect 44132 -15549 48334 -15473
rect 44098 -15575 48368 -15549
rect 44098 -15609 44158 -15575
rect 48308 -15609 48368 -15575
<< viali >>
rect 46637 -14504 47854 -14467
rect 44500 -15352 45707 -15345
rect 45707 -15352 45865 -15345
rect 45865 -15352 46291 -15345
rect 46291 -15352 46363 -15345
rect 44500 -15380 46363 -15352
rect 46616 -15401 48018 -15355
<< metal1 >>
rect 44011 -14426 48071 -14409
rect 44011 -14543 45331 -14426
rect 45670 -14467 48071 -14426
rect 45670 -14504 46637 -14467
rect 47854 -14504 48071 -14467
rect 45670 -14543 48071 -14504
rect 44011 -14555 48071 -14543
rect 44011 -15325 46402 -15311
rect 44011 -15345 44729 -15325
rect 45070 -15345 46402 -15325
rect 44011 -15380 44500 -15345
rect 46363 -15380 46402 -15345
rect 44011 -15444 44729 -15380
rect 45070 -15444 46402 -15380
rect 44011 -15457 46402 -15444
rect 46594 -15355 48070 -15311
rect 46594 -15401 46616 -15355
rect 48018 -15401 48070 -15355
rect 46594 -15457 48070 -15401
<< via1 >>
rect 45331 -14543 45670 -14426
rect 44729 -15345 45070 -15325
rect 44729 -15380 45070 -15345
rect 44729 -15444 45070 -15380
<< metal2 >>
rect 45285 -14336 45685 -14318
rect 45285 -14543 45302 -14336
rect 45670 -14543 45685 -14336
rect 45285 -14555 45685 -14543
rect 44685 -15325 45085 -15311
rect 44685 -15512 44701 -15325
rect 45070 -15512 45085 -15325
rect 44685 -15525 45085 -15512
rect 46485 -15673 46885 -15655
rect 46485 -15935 46506 -15673
rect 46868 -15935 46885 -15673
rect 46485 -15952 46885 -15935
<< via2 >>
rect 45302 -14426 45670 -14336
rect 45302 -14543 45331 -14426
rect 45331 -14543 45670 -14426
rect 44701 -15444 44729 -15325
rect 44729 -15444 45070 -15325
rect 44701 -15512 45070 -15444
rect 46506 -15935 46868 -15673
<< metal3 >>
rect 45285 -14336 45685 -14318
rect 45285 -14543 45302 -14336
rect 45670 -14543 45685 -14336
rect 45285 -14555 45685 -14543
rect 44685 -15325 45085 -15311
rect 44685 -15512 44701 -15325
rect 45070 -15512 45085 -15325
rect 44685 -15525 45085 -15512
rect 46485 -15673 46885 -15655
rect 46485 -15935 46506 -15673
rect 46868 -15935 46885 -15673
rect 46485 -15952 46885 -15935
<< labels >>
flabel metal1 44011 -14555 44167 -14409 0 FreeSans 800 0 0 0 avss
port 5 nsew
flabel metal1 44011 -15457 44167 -15311 0 FreeSans 800 0 0 0 avdd
port 4 nsew
<< end >>
