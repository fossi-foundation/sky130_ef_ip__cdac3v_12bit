magic
tech sky130A
magscale 1 2
timestamp 1747669346
<< locali >>
rect 54594 16058 54867 16072
rect 54594 15958 54614 16058
rect 54849 15958 54867 16058
rect 57090 16058 57363 16072
rect 54594 15938 54867 15958
rect 57090 15958 57110 16058
rect 57345 15958 57363 16058
rect 59586 16058 59859 16072
rect 57090 15938 57363 15958
rect 59586 15958 59606 16058
rect 59841 15958 59859 16058
rect 62082 16058 62355 16072
rect 59586 15938 59859 15958
rect 62082 15958 62102 16058
rect 62337 15958 62355 16058
rect 64578 16058 64851 16072
rect 62082 15938 62355 15958
rect 64578 15958 64598 16058
rect 64833 15958 64851 16058
rect 67074 16058 67347 16072
rect 64578 15938 64851 15958
rect 67074 15958 67094 16058
rect 67329 15958 67347 16058
rect 69570 16058 69843 16072
rect 67074 15938 67347 15958
rect 69570 15958 69590 16058
rect 69825 15958 69843 16058
rect 72066 16058 72339 16072
rect 69570 15938 69843 15958
rect 72066 15958 72086 16058
rect 72321 15958 72339 16058
rect 74562 16058 74835 16072
rect 72066 15938 72339 15958
rect 74562 15958 74582 16058
rect 74817 15958 74835 16058
rect 77058 16058 77331 16072
rect 74562 15938 74835 15958
rect 77058 15958 77078 16058
rect 77313 15958 77331 16058
rect 79554 16058 79827 16072
rect 77058 15938 77331 15958
rect 79554 15958 79574 16058
rect 79809 15958 79827 16058
rect 82050 16058 82323 16072
rect 79554 15938 79827 15958
rect 82050 15958 82070 16058
rect 82305 15958 82323 16058
rect 84546 16058 84819 16072
rect 82050 15938 82323 15958
rect 84546 15958 84566 16058
rect 84801 15958 84819 16058
rect 87042 16058 87315 16072
rect 84546 15938 84819 15958
rect 87042 15958 87062 16058
rect 87297 15958 87315 16058
rect 87042 15938 87315 15958
rect 56410 15240 56532 15252
rect 54387 15148 54649 15162
rect 54010 15132 54075 15144
rect 54010 14926 54017 15132
rect 54068 14926 54075 15132
rect 54387 15127 54407 15148
rect 54343 15060 54407 15127
rect 54387 15048 54407 15060
rect 54632 15048 54649 15148
rect 56410 15074 56420 15240
rect 56521 15074 56532 15240
rect 56410 15062 56532 15074
rect 58906 15240 59028 15252
rect 58906 15074 58916 15240
rect 59017 15074 59028 15240
rect 58906 15062 59028 15074
rect 61402 15240 61524 15252
rect 61402 15074 61412 15240
rect 61513 15074 61524 15240
rect 61402 15062 61524 15074
rect 63898 15240 64020 15252
rect 63898 15074 63908 15240
rect 64009 15074 64020 15240
rect 63898 15062 64020 15074
rect 66394 15240 66516 15252
rect 66394 15074 66404 15240
rect 66505 15074 66516 15240
rect 66394 15062 66516 15074
rect 68890 15240 69012 15252
rect 68890 15074 68900 15240
rect 69001 15074 69012 15240
rect 68890 15062 69012 15074
rect 71386 15240 71508 15252
rect 71386 15074 71396 15240
rect 71497 15074 71508 15240
rect 71386 15062 71508 15074
rect 73882 15240 74004 15252
rect 73882 15074 73892 15240
rect 73993 15074 74004 15240
rect 73882 15062 74004 15074
rect 76378 15240 76500 15252
rect 76378 15074 76388 15240
rect 76489 15074 76500 15240
rect 76378 15062 76500 15074
rect 78874 15240 78996 15252
rect 78874 15074 78884 15240
rect 78985 15074 78996 15240
rect 78874 15062 78996 15074
rect 81370 15240 81492 15252
rect 81370 15074 81380 15240
rect 81481 15074 81492 15240
rect 81370 15062 81492 15074
rect 83866 15240 83988 15252
rect 83866 15074 83876 15240
rect 83977 15074 83988 15240
rect 83866 15062 83988 15074
rect 86362 15240 86484 15252
rect 86362 15074 86372 15240
rect 86473 15074 86484 15240
rect 86362 15062 86484 15074
rect 88858 15240 88980 15252
rect 88858 15074 88868 15240
rect 88969 15074 88980 15240
rect 88858 15062 88980 15074
rect 54387 15028 54649 15048
rect 54010 14914 54075 14926
<< viali >>
rect 54614 15958 54849 16058
rect 56535 15873 56611 16049
rect 57110 15958 57345 16058
rect 59031 15873 59107 16049
rect 59606 15958 59841 16058
rect 61527 15873 61603 16049
rect 62102 15958 62337 16058
rect 64023 15873 64099 16049
rect 64598 15958 64833 16058
rect 66519 15873 66595 16049
rect 67094 15958 67329 16058
rect 69015 15873 69091 16049
rect 69590 15958 69825 16058
rect 71511 15873 71587 16049
rect 72086 15958 72321 16058
rect 74007 15873 74083 16049
rect 74582 15958 74817 16058
rect 76503 15873 76579 16049
rect 77078 15958 77313 16058
rect 78999 15873 79075 16049
rect 79574 15958 79809 16058
rect 81495 15873 81571 16049
rect 82070 15958 82305 16058
rect 83991 15873 84067 16049
rect 84566 15958 84801 16058
rect 86487 15873 86563 16049
rect 87062 15958 87297 16058
rect 88983 15873 89059 16049
rect 54017 14926 54068 15132
rect 54407 15048 54632 15148
rect 56420 15074 56521 15240
rect 58916 15074 59017 15240
rect 61412 15074 61513 15240
rect 63908 15074 64009 15240
rect 66404 15074 66505 15240
rect 68900 15074 69001 15240
rect 71396 15074 71497 15240
rect 73892 15074 73993 15240
rect 76388 15074 76489 15240
rect 78884 15074 78985 15240
rect 81380 15074 81481 15240
rect 83876 15074 83977 15240
rect 86372 15074 86473 15240
rect 88868 15074 88969 15240
<< metal1 >>
rect 53884 16253 56852 16401
rect 57019 16253 59348 16401
rect 59515 16253 61844 16401
rect 62011 16253 64340 16401
rect 64507 16253 66836 16401
rect 67003 16253 69332 16401
rect 69499 16253 71828 16401
rect 71995 16253 74324 16401
rect 74491 16253 76820 16401
rect 76987 16253 79316 16401
rect 79483 16253 81812 16401
rect 81979 16253 84308 16401
rect 84475 16253 86804 16401
rect 86971 16253 89312 16401
rect 54594 16058 54867 16072
rect 54594 15958 54614 16058
rect 54849 16038 54867 16058
rect 56520 16049 56628 16070
rect 56520 16038 56535 16049
rect 54849 15981 56535 16038
rect 54849 15958 54867 15981
rect 54594 15938 54867 15958
rect 56520 15873 56535 15981
rect 56611 15873 56628 16049
rect 57090 16058 57363 16072
rect 57090 15958 57110 16058
rect 57345 16038 57363 16058
rect 59016 16049 59124 16070
rect 59016 16038 59031 16049
rect 57345 15981 59031 16038
rect 57345 15958 57363 15981
rect 57090 15938 57363 15958
rect 54369 15790 54516 15865
rect 56520 15855 56628 15873
rect 59016 15873 59031 15981
rect 59107 15873 59124 16049
rect 59586 16058 59859 16072
rect 59586 15958 59606 16058
rect 59841 16038 59859 16058
rect 61512 16049 61620 16070
rect 61512 16038 61527 16049
rect 59841 15981 61527 16038
rect 59841 15958 59859 15981
rect 59586 15938 59859 15958
rect 59016 15855 59124 15873
rect 61512 15873 61527 15981
rect 61603 15873 61620 16049
rect 62082 16058 62355 16072
rect 62082 15958 62102 16058
rect 62337 16038 62355 16058
rect 64008 16049 64116 16070
rect 64008 16038 64023 16049
rect 62337 15981 64023 16038
rect 62337 15958 62355 15981
rect 62082 15938 62355 15958
rect 61512 15855 61620 15873
rect 64008 15873 64023 15981
rect 64099 15873 64116 16049
rect 64578 16058 64851 16072
rect 64578 15958 64598 16058
rect 64833 16038 64851 16058
rect 66504 16049 66612 16070
rect 66504 16038 66519 16049
rect 64833 15981 66519 16038
rect 64833 15958 64851 15981
rect 64578 15938 64851 15958
rect 64008 15855 64116 15873
rect 66504 15873 66519 15981
rect 66595 15873 66612 16049
rect 67074 16058 67347 16072
rect 67074 15958 67094 16058
rect 67329 16038 67347 16058
rect 69000 16049 69108 16070
rect 69000 16038 69015 16049
rect 67329 15981 69015 16038
rect 67329 15958 67347 15981
rect 67074 15938 67347 15958
rect 66504 15855 66612 15873
rect 69000 15873 69015 15981
rect 69091 15873 69108 16049
rect 69570 16058 69843 16072
rect 69570 15958 69590 16058
rect 69825 16038 69843 16058
rect 71496 16049 71604 16070
rect 71496 16038 71511 16049
rect 69825 15981 71511 16038
rect 69825 15958 69843 15981
rect 69570 15938 69843 15958
rect 69000 15855 69108 15873
rect 71496 15873 71511 15981
rect 71587 15873 71604 16049
rect 72066 16058 72339 16072
rect 72066 15958 72086 16058
rect 72321 16038 72339 16058
rect 73992 16049 74100 16070
rect 73992 16038 74007 16049
rect 72321 15981 74007 16038
rect 72321 15958 72339 15981
rect 72066 15938 72339 15958
rect 71496 15855 71604 15873
rect 73992 15873 74007 15981
rect 74083 15873 74100 16049
rect 74562 16058 74835 16072
rect 74562 15958 74582 16058
rect 74817 16038 74835 16058
rect 76488 16049 76596 16070
rect 76488 16038 76503 16049
rect 74817 15981 76503 16038
rect 74817 15958 74835 15981
rect 74562 15938 74835 15958
rect 73992 15855 74100 15873
rect 76488 15873 76503 15981
rect 76579 15873 76596 16049
rect 77058 16058 77331 16072
rect 77058 15958 77078 16058
rect 77313 16038 77331 16058
rect 78984 16049 79092 16070
rect 78984 16038 78999 16049
rect 77313 15981 78999 16038
rect 77313 15958 77331 15981
rect 77058 15938 77331 15958
rect 76488 15855 76596 15873
rect 78984 15873 78999 15981
rect 79075 15873 79092 16049
rect 79554 16058 79827 16072
rect 79554 15958 79574 16058
rect 79809 16038 79827 16058
rect 81480 16049 81588 16070
rect 81480 16038 81495 16049
rect 79809 15981 81495 16038
rect 79809 15958 79827 15981
rect 79554 15938 79827 15958
rect 78984 15855 79092 15873
rect 81480 15873 81495 15981
rect 81571 15873 81588 16049
rect 82050 16058 82323 16072
rect 82050 15958 82070 16058
rect 82305 16038 82323 16058
rect 83976 16049 84084 16070
rect 83976 16038 83991 16049
rect 82305 15981 83991 16038
rect 82305 15958 82323 15981
rect 82050 15938 82323 15958
rect 81480 15855 81588 15873
rect 83976 15873 83991 15981
rect 84067 15873 84084 16049
rect 84546 16058 84819 16072
rect 84546 15958 84566 16058
rect 84801 16038 84819 16058
rect 86472 16049 86580 16070
rect 86472 16038 86487 16049
rect 84801 15981 86487 16038
rect 84801 15958 84819 15981
rect 84546 15938 84819 15958
rect 83976 15855 84084 15873
rect 86472 15873 86487 15981
rect 86563 15873 86580 16049
rect 87042 16058 87315 16072
rect 87042 15958 87062 16058
rect 87297 16038 87315 16058
rect 88968 16049 89076 16070
rect 88968 16038 88983 16049
rect 87297 15981 88983 16038
rect 87297 15958 87315 15981
rect 87042 15938 87315 15958
rect 86472 15855 86580 15873
rect 88968 15873 88983 15981
rect 89059 15873 89076 16049
rect 88968 15855 89076 15873
rect 53886 15717 89314 15790
rect 53885 15439 89312 15689
rect 56410 15240 56532 15252
rect 54387 15148 54649 15162
rect 54010 15133 54075 15144
rect 54010 14926 54011 15133
rect 54387 15048 54407 15148
rect 54632 15131 54649 15148
rect 56410 15131 56420 15240
rect 54632 15087 56420 15131
rect 54632 15048 54649 15087
rect 56410 15074 56420 15087
rect 56521 15074 56532 15240
rect 56410 15062 56532 15074
rect 58906 15240 59028 15252
rect 58906 15074 58916 15240
rect 59017 15074 59028 15240
rect 58906 15062 59028 15074
rect 61402 15240 61524 15252
rect 61402 15074 61412 15240
rect 61513 15074 61524 15240
rect 61402 15062 61524 15074
rect 63898 15240 64020 15252
rect 63898 15074 63908 15240
rect 64009 15074 64020 15240
rect 63898 15062 64020 15074
rect 66394 15240 66516 15252
rect 66394 15074 66404 15240
rect 66505 15074 66516 15240
rect 66394 15062 66516 15074
rect 68890 15240 69012 15252
rect 68890 15074 68900 15240
rect 69001 15074 69012 15240
rect 68890 15062 69012 15074
rect 71386 15240 71508 15252
rect 71386 15074 71396 15240
rect 71497 15074 71508 15240
rect 71386 15062 71508 15074
rect 73882 15240 74004 15252
rect 73882 15074 73892 15240
rect 73993 15074 74004 15240
rect 73882 15062 74004 15074
rect 76378 15240 76500 15252
rect 76378 15074 76388 15240
rect 76489 15074 76500 15240
rect 76378 15062 76500 15074
rect 78874 15240 78996 15252
rect 78874 15074 78884 15240
rect 78985 15074 78996 15240
rect 78874 15062 78996 15074
rect 81370 15240 81492 15252
rect 81370 15074 81380 15240
rect 81481 15074 81492 15240
rect 81370 15062 81492 15074
rect 83866 15240 83988 15252
rect 83866 15074 83876 15240
rect 83977 15074 83988 15240
rect 83866 15062 83988 15074
rect 86362 15240 86484 15252
rect 86362 15074 86372 15240
rect 86473 15074 86484 15240
rect 86362 15062 86484 15074
rect 88858 15240 88980 15252
rect 88858 15074 88868 15240
rect 88969 15074 88980 15240
rect 88858 15062 88980 15074
rect 54387 15028 54649 15048
rect 54010 14914 54075 14926
rect 53886 14727 56852 14875
rect 57019 14727 59348 14875
rect 59515 14727 61844 14875
rect 62011 14727 64340 14875
rect 64507 14727 66836 14875
rect 67003 14727 69332 14875
rect 69499 14727 71828 14875
rect 71995 14727 74324 14875
rect 74491 14727 76820 14875
rect 76987 14727 79316 14875
rect 79483 14727 81812 14875
rect 81979 14727 84308 14875
rect 84475 14727 86804 14875
rect 86971 14727 89312 14875
<< via1 >>
rect 56852 16253 57019 16401
rect 59348 16253 59515 16401
rect 61844 16253 62011 16401
rect 64340 16253 64507 16401
rect 66836 16253 67003 16401
rect 69332 16253 69499 16401
rect 71828 16253 71995 16401
rect 74324 16253 74491 16401
rect 76820 16253 76987 16401
rect 79316 16253 79483 16401
rect 81812 16253 81979 16401
rect 84308 16253 84475 16401
rect 86804 16253 86971 16401
rect 54614 15958 54849 16058
rect 57110 15958 57345 16058
rect 59606 15958 59841 16058
rect 62102 15958 62337 16058
rect 64598 15958 64833 16058
rect 67094 15958 67329 16058
rect 69590 15958 69825 16058
rect 72086 15958 72321 16058
rect 74582 15958 74817 16058
rect 77078 15958 77313 16058
rect 79574 15958 79809 16058
rect 82070 15958 82305 16058
rect 84566 15958 84801 16058
rect 87062 15958 87297 16058
rect 54011 15132 54075 15133
rect 54011 14926 54017 15132
rect 54017 14926 54068 15132
rect 54068 14926 54075 15132
rect 56420 15074 56521 15240
rect 58916 15074 59017 15240
rect 61412 15074 61513 15240
rect 63908 15074 64009 15240
rect 66404 15074 66505 15240
rect 68900 15074 69001 15240
rect 71396 15074 71497 15240
rect 73892 15074 73993 15240
rect 76388 15074 76489 15240
rect 78884 15074 78985 15240
rect 81380 15074 81481 15240
rect 83876 15074 83977 15240
rect 86372 15074 86473 15240
rect 88868 15074 88969 15240
rect 56852 14727 57019 14875
rect 59348 14727 59515 14875
rect 61844 14727 62011 14875
rect 64340 14727 64507 14875
rect 66836 14727 67003 14875
rect 69332 14727 69499 14875
rect 71828 14727 71995 14875
rect 74324 14727 74491 14875
rect 76820 14727 76987 14875
rect 79316 14727 79483 14875
rect 81812 14727 81979 14875
rect 84308 14727 84475 14875
rect 86804 14727 86971 14875
<< metal2 >>
rect 54711 16073 54755 16424
rect 56852 16401 57019 16412
rect 54594 16058 54866 16073
rect 54594 15958 54614 16058
rect 54849 15958 54866 16058
rect 54594 15938 54866 15958
rect 56410 15240 56532 15252
rect 54010 15133 54075 15144
rect 54010 14926 54011 15133
rect 56410 15074 56420 15240
rect 56521 15074 56532 15240
rect 56410 15062 56532 15074
rect 54010 14914 54075 14926
rect 54021 14707 54062 14914
rect 56450 14704 56494 15062
rect 56852 14875 57019 16253
rect 57207 16073 57251 16424
rect 59348 16401 59515 16412
rect 57090 16058 57362 16073
rect 57090 15958 57110 16058
rect 57345 15958 57362 16058
rect 57090 15938 57362 15958
rect 58906 15240 59028 15252
rect 58906 15074 58916 15240
rect 59017 15074 59028 15240
rect 58906 15062 59028 15074
rect 56852 14719 57019 14727
rect 58946 14704 58990 15062
rect 59348 14875 59515 16253
rect 59703 16073 59747 16424
rect 61844 16401 62011 16412
rect 59586 16058 59858 16073
rect 59586 15958 59606 16058
rect 59841 15958 59858 16058
rect 59586 15938 59858 15958
rect 61402 15240 61524 15252
rect 61402 15074 61412 15240
rect 61513 15074 61524 15240
rect 61402 15062 61524 15074
rect 59348 14719 59515 14727
rect 61442 14704 61486 15062
rect 61844 14875 62011 16253
rect 62199 16073 62243 16424
rect 64340 16401 64507 16412
rect 62082 16058 62354 16073
rect 62082 15958 62102 16058
rect 62337 15958 62354 16058
rect 62082 15938 62354 15958
rect 63898 15240 64020 15252
rect 63898 15074 63908 15240
rect 64009 15074 64020 15240
rect 63898 15062 64020 15074
rect 61844 14719 62011 14727
rect 63938 14704 63982 15062
rect 64340 14875 64507 16253
rect 64695 16073 64739 16424
rect 66836 16401 67003 16412
rect 64578 16058 64850 16073
rect 64578 15958 64598 16058
rect 64833 15958 64850 16058
rect 64578 15938 64850 15958
rect 66394 15240 66516 15252
rect 66394 15074 66404 15240
rect 66505 15074 66516 15240
rect 66394 15062 66516 15074
rect 64340 14719 64507 14727
rect 66434 14704 66478 15062
rect 66836 14875 67003 16253
rect 67191 16073 67235 16424
rect 69332 16401 69499 16412
rect 67074 16058 67346 16073
rect 67074 15958 67094 16058
rect 67329 15958 67346 16058
rect 67074 15938 67346 15958
rect 68890 15240 69012 15252
rect 68890 15074 68900 15240
rect 69001 15074 69012 15240
rect 68890 15062 69012 15074
rect 66836 14719 67003 14727
rect 68930 14704 68974 15062
rect 69332 14875 69499 16253
rect 69687 16073 69731 16424
rect 71828 16401 71995 16412
rect 69570 16058 69842 16073
rect 69570 15958 69590 16058
rect 69825 15958 69842 16058
rect 69570 15938 69842 15958
rect 71386 15240 71508 15252
rect 71386 15074 71396 15240
rect 71497 15074 71508 15240
rect 71386 15062 71508 15074
rect 69332 14719 69499 14727
rect 71426 14704 71470 15062
rect 71828 14875 71995 16253
rect 72183 16073 72227 16424
rect 74324 16401 74491 16412
rect 72066 16058 72338 16073
rect 72066 15958 72086 16058
rect 72321 15958 72338 16058
rect 72066 15938 72338 15958
rect 73882 15240 74004 15252
rect 73882 15074 73892 15240
rect 73993 15074 74004 15240
rect 73882 15062 74004 15074
rect 71828 14719 71995 14727
rect 73922 14704 73966 15062
rect 74324 14875 74491 16253
rect 74679 16073 74723 16424
rect 76820 16401 76987 16412
rect 74562 16058 74834 16073
rect 74562 15958 74582 16058
rect 74817 15958 74834 16058
rect 74562 15938 74834 15958
rect 76378 15240 76500 15252
rect 76378 15074 76388 15240
rect 76489 15074 76500 15240
rect 76378 15062 76500 15074
rect 74324 14719 74491 14727
rect 76418 14704 76462 15062
rect 76820 14875 76987 16253
rect 77175 16073 77219 16424
rect 79316 16401 79483 16412
rect 77058 16058 77330 16073
rect 77058 15958 77078 16058
rect 77313 15958 77330 16058
rect 77058 15938 77330 15958
rect 78874 15240 78996 15252
rect 78874 15074 78884 15240
rect 78985 15074 78996 15240
rect 78874 15062 78996 15074
rect 76820 14719 76987 14727
rect 78914 14704 78958 15062
rect 79316 14875 79483 16253
rect 79671 16073 79715 16424
rect 81812 16401 81979 16412
rect 79554 16058 79826 16073
rect 79554 15958 79574 16058
rect 79809 15958 79826 16058
rect 79554 15938 79826 15958
rect 81370 15240 81492 15252
rect 81370 15074 81380 15240
rect 81481 15074 81492 15240
rect 81370 15062 81492 15074
rect 79316 14719 79483 14727
rect 81410 14704 81454 15062
rect 81812 14875 81979 16253
rect 82167 16073 82211 16424
rect 84308 16401 84475 16412
rect 82050 16058 82322 16073
rect 82050 15958 82070 16058
rect 82305 15958 82322 16058
rect 82050 15938 82322 15958
rect 83866 15240 83988 15252
rect 83866 15074 83876 15240
rect 83977 15074 83988 15240
rect 83866 15062 83988 15074
rect 81812 14719 81979 14727
rect 83906 14704 83950 15062
rect 84308 14875 84475 16253
rect 84663 16073 84707 16424
rect 86804 16401 86971 16412
rect 84546 16058 84818 16073
rect 84546 15958 84566 16058
rect 84801 15958 84818 16058
rect 84546 15938 84818 15958
rect 86362 15240 86484 15252
rect 86362 15074 86372 15240
rect 86473 15074 86484 15240
rect 86362 15062 86484 15074
rect 84308 14719 84475 14727
rect 86402 14704 86446 15062
rect 86804 14875 86971 16253
rect 87159 16073 87203 16424
rect 87042 16058 87314 16073
rect 87042 15958 87062 16058
rect 87297 15958 87314 16058
rect 87042 15938 87314 15958
rect 88858 15240 88980 15252
rect 88858 15074 88868 15240
rect 88969 15074 88980 15240
rect 88858 15062 88980 15074
rect 86804 14719 86971 14727
rect 88898 14704 88942 15062
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 1 0 63968 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_1
timestamp 1747669346
transform 1 0 56480 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_2
timestamp 1747669346
transform 1 0 58976 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_3
timestamp 1747669346
transform 1 0 61472 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_4
timestamp 1747669346
transform 1 0 66464 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_5
timestamp 1747669346
transform 1 0 68960 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_6
timestamp 1747669346
transform 1 0 71456 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_7
timestamp 1747669346
transform 1 0 78944 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_8
timestamp 1747669346
transform 1 0 73952 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_9
timestamp 1747669346
transform 1 0 76448 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_10
timestamp 1747669346
transform 1 0 81440 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_11
timestamp 1747669346
transform 1 0 86432 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_12
timestamp 1747669346
transform 1 0 83936 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_13
timestamp 1747669346
transform 1 0 88928 0 1 14750
box -66 -43 450 897
use sky130_fd_sc_hvl__decap_4  sky130_fd_sc_hvl__decap_4_14
timestamp 1747669346
transform 1 0 53984 0 -1 16378
box -66 -43 450 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 1 0 63968 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_1
timestamp 1747669346
transform 1 0 56480 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_2
timestamp 1747669346
transform 1 0 58976 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_3
timestamp 1747669346
transform 1 0 61472 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_4
timestamp 1747669346
transform 1 0 66464 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_5
timestamp 1747669346
transform 1 0 68960 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_6
timestamp 1747669346
transform 1 0 71456 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_7
timestamp 1747669346
transform 1 0 78944 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_8
timestamp 1747669346
transform 1 0 73952 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_9
timestamp 1747669346
transform 1 0 76448 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_10
timestamp 1747669346
transform 1 0 81440 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_11
timestamp 1747669346
transform 1 0 86432 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_12
timestamp 1747669346
transform 1 0 83936 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__diode_2  sky130_fd_sc_hvl__diode_2_13
timestamp 1747669346
transform 1 0 88928 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_1  sky130_fd_sc_hvl__fill_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 1 0 53888 0 -1 16378
box -66 -43 162 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 1 0 64160 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_1
timestamp 1747669346
transform 1 0 56672 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_2
timestamp 1747669346
transform 1 0 59168 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_3
timestamp 1747669346
transform 1 0 61664 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_4
timestamp 1747669346
transform 1 0 66656 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_5
timestamp 1747669346
transform 1 0 69152 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_6
timestamp 1747669346
transform 1 0 71648 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_7
timestamp 1747669346
transform 1 0 76640 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_8
timestamp 1747669346
transform 1 0 74144 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_9
timestamp 1747669346
transform 1 0 81632 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_10
timestamp 1747669346
transform 1 0 79136 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_11
timestamp 1747669346
transform 1 0 89120 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_12
timestamp 1747669346
transform 1 0 84128 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__fill_2  sky130_fd_sc_hvl__fill_2_13
timestamp 1747669346
transform 1 0 86624 0 -1 16378
box -66 -43 258 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform -1 0 54368 0 1 14750
box -66 -43 546 897
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 1 0 59360 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_1
timestamp 1747669346
transform 1 0 54368 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_2
timestamp 1747669346
transform 1 0 56864 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_3
timestamp 1747669346
transform 1 0 64352 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_4
timestamp 1747669346
transform 1 0 61856 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_5
timestamp 1747669346
transform 1 0 66848 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_6
timestamp 1747669346
transform 1 0 69344 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_7
timestamp 1747669346
transform 1 0 71840 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_8
timestamp 1747669346
transform 1 0 74336 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_9
timestamp 1747669346
transform 1 0 76832 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_10
timestamp 1747669346
transform 1 0 81824 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_11
timestamp 1747669346
transform 1 0 79328 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_12
timestamp 1747669346
transform 1 0 84320 0 -1 16378
box -66 -43 2178 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_13
timestamp 1747669346
transform 1 0 86816 0 -1 16378
box -66 -43 2178 1671
<< labels >>
flabel metal2 54711 16289 54755 16424 0 FreeSans 480 90 0 0 HOLD
port 0 nsew
flabel metal2 57207 16289 57251 16424 0 FreeSans 480 90 0 0 RST
port 1 nsew
flabel metal2 59703 16289 59747 16424 0 FreeSans 480 90 0 0 SEL0
port 2 nsew
flabel metal2 62199 16289 62243 16424 0 FreeSans 480 90 0 0 SEL1
port 3 nsew
flabel metal2 64695 16289 64739 16424 0 FreeSans 480 90 0 0 SEL2
port 4 nsew
flabel metal2 67191 16289 67235 16424 0 FreeSans 480 90 0 0 SEL3
port 5 nsew
flabel metal2 69687 16289 69731 16424 0 FreeSans 480 90 0 0 SEL4
port 6 nsew
flabel metal2 72183 16289 72227 16424 0 FreeSans 480 90 0 0 SEL5
port 7 nsew
flabel metal2 74679 16289 74723 16424 0 FreeSans 480 90 0 0 SEL6
port 8 nsew
flabel metal2 77175 16289 77219 16424 0 FreeSans 480 90 0 0 SEL7
port 9 nsew
flabel metal2 79671 16289 79715 16424 0 FreeSans 480 90 0 0 SEL8
port 10 nsew
flabel metal2 82167 16289 82211 16424 0 FreeSans 480 90 0 0 SEL9
port 11 nsew
flabel metal2 84663 16289 84707 16424 0 FreeSans 480 90 0 0 SEL10
port 12 nsew
flabel metal2 87159 16289 87203 16424 0 FreeSans 480 90 0 0 SEL11
port 13 nsew
flabel metal2 56450 14704 56494 14839 0 FreeSans 480 90 0 0 HOLD_3P3
port 14 nsew
flabel metal2 58946 14704 58990 14839 0 FreeSans 480 90 0 0 RST_3P3
port 15 nsew
flabel metal2 61442 14704 61486 14839 0 FreeSans 480 90 0 0 SEL0_3P3
port 16 nsew
flabel metal2 63938 14704 63982 14839 0 FreeSans 480 90 0 0 SEL1_3P3
port 17 nsew
flabel metal2 66434 14704 66478 14839 0 FreeSans 480 90 0 0 SEL2_3P3
port 18 nsew
flabel metal2 68930 14704 68974 14839 0 FreeSans 480 90 0 0 SEL3_3P3
port 19 nsew
flabel metal2 71426 14704 71470 14839 0 FreeSans 480 90 0 0 SEL4_3P3
port 20 nsew
flabel metal2 73922 14704 73966 14839 0 FreeSans 480 90 0 0 SEL5_3P3
port 21 nsew
flabel metal2 76418 14704 76462 14839 0 FreeSans 480 90 0 0 SEL6_3P3
port 22 nsew
flabel metal2 78914 14704 78958 14839 0 FreeSans 480 90 0 0 SEL7_3P3
port 23 nsew
flabel metal2 81410 14704 81454 14839 0 FreeSans 480 90 0 0 SEL8_3P3
port 24 nsew
flabel metal2 83906 14704 83950 14839 0 FreeSans 480 90 0 0 SEL9_3P3
port 25 nsew
flabel metal2 88898 14704 88942 14839 0 FreeSans 480 90 0 0 SEL11_3P3
port 27 nsew
flabel metal1 54368 14727 54515 14875 0 FreeSans 480 0 0 0 VSS
port 30 nsew
flabel metal1 54367 15492 54514 15640 0 FreeSans 480 0 0 0 VDD3P3
port 31 nsew
flabel metal1 54369 15717 54516 15865 0 FreeSans 480 0 0 0 VDD1P8
port 32 nsew
flabel metal2 54021 14707 54062 14862 0 FreeSans 480 90 0 0 HOLDB_3P3
port 33 nsew
flabel metal2 86404 14704 86446 14839 0 FreeSans 480 90 0 0 SEL10_3P3
port 26 nsew
<< properties >>
string MASKHINTS_HVI 53836 16421 89349 16462
<< end >>
