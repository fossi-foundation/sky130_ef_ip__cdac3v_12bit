magic
tech sky130A
magscale 1 2
timestamp 1747669346
<< error_s >>
rect 1008 -1548 4421 -1475
rect 1008 -8839 4421 -8763
<< dnwell >>
rect 1088 -1897 4341 -1555
rect 1088 -4220 4341 -3572
rect 2183 -6098 2639 -5858
rect 1088 -6506 4341 -6098
rect 1088 -8759 4341 -8411
<< nwell >>
rect 980 -1788 4451 -1548
rect 2188 -1988 2644 -1788
rect 980 -4095 4450 -3656
rect 2183 -6194 2639 -5954
rect 980 -6393 4450 -6194
rect 2180 -8514 2636 -8234
rect 979 -8763 4450 -8514
<< locali >>
rect 5183 -3949 5249 -3866
rect 5190 -4852 5239 -4840
<< viali >>
rect 5049 -3600 5228 -3558
rect 5169 -3987 5350 -3949
rect 5227 -4094 5296 -4039
rect 5238 -4358 5281 -4153
rect 5043 -4562 5222 -4520
rect 5190 -4840 5239 -4665
rect 5190 -5083 5239 -4896
rect 5043 -5228 5222 -5186
rect 5190 -5571 5239 -5384
rect 5043 -5716 5222 -5674
rect 5043 -6002 5222 -5960
rect 5190 -6292 5239 -6105
rect 5238 -6562 5281 -6357
rect 5227 -6676 5296 -6623
rect 5169 -6766 5350 -6728
<< metal1 >>
rect 4488 -1642 4540 -1631
rect 2778 -1732 4488 -1696
rect 2780 -1816 2816 -1732
rect 4488 -1794 4540 -1781
rect 4488 -1844 4540 -1833
rect 2898 -1947 4488 -1904
rect 4488 -1996 4540 -1983
rect 4480 -3941 4532 -3930
rect 2769 -4027 4480 -3990
rect 2769 -4113 2806 -4027
rect 4480 -4093 4532 -4080
rect 4479 -4141 4531 -4130
rect 2883 -4259 4479 -4222
rect 4479 -4293 4531 -4280
rect 4492 -6175 4545 -6167
rect 2770 -6311 4492 -6279
rect 4544 -6311 4545 -6175
rect 2770 -6319 4545 -6311
rect 2770 -6400 2810 -6319
rect 4492 -6321 4545 -6319
rect 2900 -6384 4545 -6376
rect 2900 -6416 4492 -6384
rect 4544 -6520 4545 -6384
rect 4492 -6530 4545 -6520
rect 4846 -8501 4997 -1545
rect 5405 -1625 5469 -1552
rect 5182 -1703 5234 -1692
rect 5399 -1825 5475 -1625
rect 5182 -1855 5234 -1842
rect 5285 -1844 5337 -1833
rect 5191 -3548 5228 -1855
rect 5285 -1996 5337 -1983
rect 5034 -3558 5242 -3548
rect 5034 -3600 5049 -3558
rect 5228 -3600 5242 -3558
rect 5034 -3608 5242 -3600
rect 5296 -3942 5334 -1996
rect 5157 -3949 5362 -3942
rect 5157 -3987 5169 -3949
rect 5350 -3987 5362 -3949
rect 5157 -3994 5362 -3987
rect 5204 -4039 5323 -4026
rect 5204 -4057 5227 -4039
rect 5112 -4094 5227 -4057
rect 5296 -4094 5323 -4039
rect 5112 -4105 5323 -4094
rect 5112 -4510 5154 -4105
rect 5227 -4153 5296 -4134
rect 5227 -4358 5238 -4153
rect 5281 -4213 5296 -4153
rect 5405 -4213 5469 -1825
rect 5281 -4276 5469 -4213
rect 5281 -4358 5296 -4276
rect 5227 -4373 5296 -4358
rect 5028 -4520 5236 -4510
rect 5028 -4562 5043 -4520
rect 5222 -4562 5236 -4520
rect 5028 -4570 5236 -4562
rect 5182 -4652 5248 -4639
rect 5165 -4764 5182 -4716
rect 5248 -4764 5347 -4716
rect 5182 -4853 5248 -4840
rect 5182 -4893 5248 -4882
rect 5182 -5096 5248 -5084
rect 5182 -5178 5248 -5177
rect 5028 -5238 5039 -5178
rect 5234 -5238 5248 -5178
rect 5182 -5384 5248 -5238
rect 5182 -5571 5190 -5384
rect 5239 -5571 5248 -5384
rect 5182 -5584 5248 -5571
rect 5028 -5726 5037 -5666
rect 5226 -5726 5236 -5666
rect 5028 -6010 5035 -5950
rect 5227 -6010 5236 -5950
rect 5182 -6105 5248 -6092
rect 5182 -6226 5190 -6105
rect 5156 -6292 5190 -6226
rect 5239 -6292 5248 -6105
rect 5156 -6306 5248 -6292
rect 5156 -6721 5193 -6306
rect 5299 -6339 5347 -4764
rect 5227 -6357 5347 -6339
rect 5227 -6562 5238 -6357
rect 5281 -6387 5347 -6357
rect 5405 -4893 5469 -4276
rect 5281 -6562 5296 -6387
rect 5227 -6581 5296 -6562
rect 5405 -6609 5469 -5084
rect 5221 -6623 5469 -6609
rect 5221 -6676 5227 -6623
rect 5296 -6676 5469 -6623
rect 5221 -6689 5469 -6676
rect 5156 -6773 5169 -6721
rect 5350 -6773 5362 -6721
rect 5156 -6777 5193 -6773
rect 4846 -8756 4997 -8725
rect 5405 -8758 5469 -6689
rect 5560 -2039 5711 -1543
rect 5560 -8756 5711 -2236
<< via1 >>
rect 4488 -1781 4540 -1642
rect 4488 -1983 4540 -1844
rect 1629 -2166 2685 -2098
rect 2970 -3620 4008 -3564
rect 4480 -4080 4532 -3941
rect 4479 -4280 4531 -4141
rect 1612 -4457 2005 -4388
rect 2970 -5880 4008 -5824
rect 4492 -6311 4544 -6175
rect 4492 -6520 4544 -6384
rect 1611 -6747 2004 -6678
rect 2970 -8190 4008 -8134
rect 5182 -1842 5234 -1703
rect 5285 -1983 5337 -1844
rect 5182 -4665 5248 -4652
rect 5182 -4840 5190 -4665
rect 5190 -4840 5239 -4665
rect 5239 -4840 5248 -4665
rect 5182 -4896 5248 -4893
rect 5182 -5083 5190 -4896
rect 5190 -5083 5239 -4896
rect 5239 -5083 5248 -4896
rect 5182 -5084 5248 -5083
rect 5039 -5186 5234 -5178
rect 5039 -5228 5043 -5186
rect 5043 -5228 5222 -5186
rect 5222 -5228 5234 -5186
rect 5039 -5238 5234 -5228
rect 5037 -5674 5226 -5666
rect 5037 -5716 5043 -5674
rect 5043 -5716 5222 -5674
rect 5222 -5716 5226 -5674
rect 5037 -5726 5226 -5716
rect 5035 -5960 5227 -5950
rect 5035 -6002 5043 -5960
rect 5043 -6002 5222 -5960
rect 5222 -6002 5227 -5960
rect 5035 -6010 5227 -6002
rect 5405 -5084 5469 -4893
rect 5169 -6728 5350 -6721
rect 5169 -6766 5350 -6728
rect 5169 -6773 5350 -6766
rect 4846 -8725 4997 -8501
rect 5560 -2236 5711 -2039
<< metal2 >>
rect 4488 -1642 4540 -1631
rect 5182 -1703 5234 -1692
rect 4540 -1732 4541 -1708
rect 4540 -1762 5182 -1732
rect 4488 -1794 4540 -1781
rect 4488 -1844 4540 -1833
rect 5182 -1855 5234 -1842
rect 5285 -1844 5337 -1833
rect 4540 -1948 5285 -1910
rect 4488 -1996 4540 -1983
rect 5285 -1996 5337 -1983
rect 1609 -2014 2010 -2002
rect 1609 -2225 1627 -2014
rect 1997 -2039 2010 -2014
rect 1997 -2098 5560 -2039
rect 2685 -2166 5560 -2098
rect 1997 -2225 5560 -2166
rect 1609 -2236 5560 -2225
rect 5711 -2236 5720 -2039
rect 4114 -2364 4449 -2361
rect 3974 -2372 4449 -2364
rect 3974 -2564 4271 -2372
rect 4147 -2784 4271 -2564
rect 4426 -2784 4449 -2372
rect 4147 -2794 4449 -2784
rect 4148 -2938 4794 -2922
rect 4148 -3338 4606 -2938
rect 4769 -3338 4794 -2938
rect 4148 -3354 4794 -3338
rect 2209 -3526 4140 -3512
rect 2209 -3752 2222 -3526
rect 2596 -3564 4140 -3526
rect 2596 -3620 2970 -3564
rect 4008 -3620 4140 -3564
rect 2596 -3673 4140 -3620
rect 2596 -3752 2610 -3673
rect 2209 -3765 2610 -3752
rect 1069 -3840 1217 -3785
rect 1069 -3881 4919 -3840
rect 1069 -3916 1217 -3881
rect 4480 -3941 4532 -3930
rect 4532 -4021 4757 -3991
rect 4480 -4093 4532 -4080
rect 4479 -4141 4531 -4130
rect 1608 -4284 2010 -4269
rect 1608 -4388 1622 -4284
rect 1996 -4388 2010 -4284
rect 4531 -4227 4641 -4192
rect 4479 -4293 4531 -4280
rect 1608 -4457 1612 -4388
rect 2005 -4457 2010 -4388
rect 1608 -4498 1622 -4457
rect 1996 -4498 2010 -4457
rect 1608 -4507 2010 -4498
rect 1051 -4664 1331 -4652
rect 1051 -5065 1067 -4664
rect 4606 -5041 4641 -4227
rect 4727 -4865 4757 -4021
rect 4878 -4725 4919 -3881
rect 5182 -4652 5248 -4639
rect 4878 -4766 5182 -4725
rect 5182 -4853 5248 -4840
rect 4727 -4895 5059 -4865
rect 1051 -5084 1331 -5065
rect 4606 -5076 4896 -5041
rect 4146 -5228 4792 -5212
rect 4146 -5628 4607 -5228
rect 4770 -5628 4792 -5228
rect 4146 -5644 4792 -5628
rect 4865 -5682 4896 -5076
rect 5022 -5178 5059 -4895
rect 5182 -4893 5248 -4881
rect 5405 -4893 5469 -4881
rect 5248 -5016 5405 -4962
rect 5182 -5096 5248 -5084
rect 5405 -5095 5469 -5084
rect 5022 -5238 5039 -5178
rect 5234 -5238 5248 -5178
rect 5028 -5682 5037 -5666
rect 4865 -5713 5037 -5682
rect 5028 -5726 5037 -5713
rect 5226 -5726 5236 -5666
rect 2209 -5786 4140 -5772
rect 2209 -6012 2222 -5786
rect 2596 -5824 4140 -5786
rect 2596 -5880 2970 -5824
rect 4008 -5880 4140 -5824
rect 2596 -5933 4140 -5880
rect 2596 -6012 2610 -5933
rect 5028 -5967 5035 -5950
rect 2209 -6025 2610 -6012
rect 4506 -5995 5035 -5967
rect 4506 -6167 4534 -5995
rect 5028 -6010 5035 -5995
rect 5227 -6010 5236 -5950
rect 4492 -6175 4545 -6167
rect 4544 -6311 4545 -6175
rect 4492 -6321 4545 -6311
rect 4492 -6384 4545 -6376
rect 4544 -6520 4545 -6384
rect 4492 -6530 4545 -6520
rect 1608 -6584 2010 -6569
rect 1608 -6678 1622 -6584
rect 1996 -6678 2010 -6584
rect 1608 -6747 1611 -6678
rect 2004 -6747 2010 -6678
rect 1608 -6798 1622 -6747
rect 1996 -6798 2010 -6747
rect 4502 -6733 4530 -6530
rect 5157 -6733 5169 -6721
rect 4502 -6761 5169 -6733
rect 5157 -6773 5169 -6761
rect 5350 -6773 5362 -6721
rect 1608 -6807 2010 -6798
rect 3911 -7358 3975 -7173
rect 3911 -7373 4111 -7358
rect 4141 -7517 4795 -7502
rect 4141 -7917 4607 -7517
rect 4770 -7917 4795 -7517
rect 4141 -7934 4795 -7917
rect 2610 -8084 4140 -8082
rect 2210 -8095 4140 -8084
rect 2210 -8298 2221 -8095
rect 2597 -8134 4140 -8095
rect 2597 -8190 2970 -8134
rect 4008 -8190 4140 -8134
rect 2597 -8243 4140 -8190
rect 2597 -8298 2610 -8243
rect 2210 -8311 2610 -8298
rect 3412 -8504 4846 -8501
rect 3409 -8520 4846 -8504
rect 3409 -8707 3426 -8520
rect 3794 -8707 4846 -8520
rect 3409 -8725 4846 -8707
rect 4997 -8725 5009 -8501
rect 3409 -8726 3810 -8725
<< via2 >>
rect 1627 -2098 1997 -2014
rect 1627 -2166 1629 -2098
rect 1629 -2166 1997 -2098
rect 1627 -2225 1997 -2166
rect 4271 -2784 4426 -2372
rect 4606 -3338 4769 -2938
rect 2222 -3752 2596 -3526
rect 1622 -4388 1996 -4284
rect 1622 -4457 1996 -4388
rect 1622 -4498 1996 -4457
rect 1067 -5065 1380 -4664
rect 4607 -5628 4770 -5228
rect 2222 -6012 2596 -5786
rect 1622 -6678 1996 -6584
rect 1622 -6747 1996 -6678
rect 1622 -6798 1996 -6747
rect 3975 -7358 4125 -6979
rect 4607 -7917 4770 -7517
rect 2221 -8298 2597 -8095
rect 3426 -8707 3794 -8520
<< metal3 >>
rect 1047 -4664 1397 -1541
rect 1047 -5065 1067 -4664
rect 1380 -5065 1397 -4664
rect 1047 -8752 1397 -5065
rect 1610 -2014 2010 -1545
rect 1610 -2225 1627 -2014
rect 1997 -2225 2010 -2014
rect 1610 -4284 2010 -2225
rect 1610 -4498 1622 -4284
rect 1996 -4498 2010 -4284
rect 1610 -6584 2010 -4498
rect 1610 -6798 1622 -6584
rect 1996 -6798 2010 -6584
rect 1610 -8757 2010 -6798
rect 2210 -3526 2610 -1545
rect 2210 -3752 2222 -3526
rect 2596 -3752 2610 -3526
rect 2210 -5786 2610 -3752
rect 2210 -6012 2222 -5786
rect 2596 -6012 2610 -5786
rect 2210 -8095 2610 -6012
rect 2210 -8298 2221 -8095
rect 2597 -8298 2610 -8095
rect 2210 -8757 2610 -8298
rect 2810 -8757 3210 -1543
rect 3410 -8520 3810 -1543
rect 3410 -8707 3426 -8520
rect 3794 -8707 3810 -8520
rect 3410 -8757 3810 -8707
rect 3959 -6979 4139 -1541
rect 3959 -7358 3975 -6979
rect 4125 -7358 4139 -6979
rect 3959 -8757 4139 -7358
rect 4259 -2372 4439 -1541
rect 4259 -2784 4271 -2372
rect 4426 -2784 4439 -2372
rect 4259 -8757 4439 -2784
rect 4591 -2938 4787 -1864
rect 4591 -3338 4606 -2938
rect 4769 -3338 4787 -2938
rect 4591 -5228 4787 -3338
rect 4591 -5628 4607 -5228
rect 4770 -5628 4787 -5228
rect 4591 -6461 4787 -5628
rect 4591 -6661 4791 -6461
rect 4591 -7517 4787 -6661
rect 4591 -7917 4607 -7517
rect 4770 -7917 4787 -7517
rect 4591 -8444 4787 -7917
use simple_analog_switch_2  simple_analog_switch_2_0 ../ip/sky130_ef_ip__analog_switches/mag
timestamp 1747669346
transform 1 0 -230 0 1 -8538
box 1210 24 4680 2176
use simple_analog_switch_2  simple_analog_switch_2_1
timestamp 1747669346
transform 1 0 -230 0 1 -3958
box 1210 24 4680 2176
use simple_analog_switch_2  simple_analog_switch_2_2
timestamp 1747669346
transform 1 0 -230 0 1 -6248
box 1210 24 4680 2176
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 0 1 4872 -1 0 -7550
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_1
timestamp 1747669346
transform 0 1 4872 -1 0 -2670
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_2
timestamp 1747669346
transform 0 1 4872 -1 0 -1902
box -66 -43 834 897
use sky130_fd_sc_hvl__decap_8  sky130_fd_sc_hvl__decap_8_3
timestamp 1747669346
transform 0 1 4872 -1 0 -6782
box -66 -43 834 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 0 1 4872 1 0 -3918
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_1
timestamp 1747669346
transform 0 1 4872 -1 0 -4878
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_2
timestamp 1747669346
transform 0 1 4872 1 0 -4878
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_3
timestamp 1747669346
transform 0 1 4872 1 0 -6318
box -66 -43 546 897
use sky130_fd_sc_hvl__inv_2  sky130_fd_sc_hvl__inv_2_5
timestamp 1747669346
transform 0 1 4872 -1 0 -5358
box -66 -43 546 897
use sky130_fd_sc_hvl__nor2_1  sky130_fd_sc_hvl__nor2_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hvl/mag
timestamp 1747669346
transform 0 1 4872 1 0 -4398
box -66 -43 546 897
use sky130_fd_sc_hvl__nor2_1  sky130_fd_sc_hvl__nor2_1_1
timestamp 1747669346
transform 0 1 4872 -1 0 -6318
box -66 -43 546 897
<< labels >>
flabel metal3 4591 -6661 4791 -6461 0 FreeSans 256 0 0 0 vo
port 2 nsew
flabel metal3 2895 -1804 3095 -1604 0 FreeSans 256 0 0 0 vdd1p8
port 1 nsew
flabel metal3 3499 -1801 3699 -1601 0 FreeSans 256 0 0 0 dvss
port 7 nsew
flabel metal3 1696 -1798 1896 -1598 0 FreeSans 256 0 0 0 vdd3p3
port 0 nsew
flabel metal3 2313 -1771 2513 -1625 0 FreeSans 256 0 0 0 vss
port 3 nsew
flabel metal3 1114 -1795 1323 -1594 0 FreeSans 480 0 0 0 cm
port 9 nsew
flabel metal3 4264 -1744 4439 -1544 0 FreeSans 256 0 0 0 b
port 5 nsew
flabel metal3 3959 -1751 4139 -1551 0 FreeSans 256 0 0 0 a
port 4 nsew
flabel metal1 5399 -1825 5475 -1625 0 FreeSans 256 90 0 0 selcm
port 8 nsew
flabel metal2 1069 -3916 1217 -3785 0 FreeSans 256 0 0 0 sel
port 6 nsew
<< end >>
