magic
tech sky130A
magscale 1 2
timestamp 1747671550
<< nwell >>
rect 1705 23500 1778 26971
rect 49417 23501 49493 26972
rect 1705 -8724 1778 -5253
rect 49417 -8725 49493 -5254
<< metal1 >>
rect 50077 23985 50242 24005
rect 50077 23492 50092 23985
rect 50229 23492 50242 23985
rect 23328 22960 23716 23111
rect 23565 22863 23716 22960
rect 27304 22954 27942 23105
rect 27304 22863 27455 22954
rect 23565 22712 27455 22863
rect 23337 22482 27875 22546
rect 23232 22240 27879 22391
rect 23243 -4144 27884 -3993
rect 23311 -4299 27900 -4235
rect 23552 -4562 27465 -4411
rect 23552 -4704 23703 -4562
rect 23371 -4855 23703 -4704
rect 27314 -4707 27465 -4562
rect 27314 -4858 27942 -4707
rect 50077 -5029 50242 23492
rect 50077 -5729 50093 -5029
rect 50228 -5729 50242 -5029
rect 50077 -5751 50242 -5729
<< via1 >>
rect 50092 23492 50229 23985
rect 50093 -5729 50228 -5029
<< metal2 >>
rect 50077 26893 50242 26919
rect 4015 26681 4215 26881
rect 11219 26683 11419 26883
rect 18424 26682 18624 26882
rect 30033 26682 30233 26882
rect 37235 26681 37435 26881
rect 44440 26680 44640 26880
rect 50077 26565 50087 26893
rect 50233 26565 50242 26893
rect 50077 23985 50242 26565
rect 50077 23492 50092 23985
rect 50229 23492 50242 23985
rect 50077 23476 50242 23492
rect 50077 -5029 50242 -5014
rect 2602 -5433 3014 -5278
rect 9806 -5433 10218 -5278
rect 15798 -5431 15988 -5281
rect 17010 -5433 17422 -5278
rect 29806 -5431 29996 -5281
rect 43022 -5436 43438 -5277
rect 7209 -5729 7588 -5579
rect 14213 -5729 14403 -5579
rect 14413 -5729 14792 -5579
rect 21217 -5729 21407 -5579
rect 21617 -5729 21996 -5579
rect 35225 -5729 35415 -5579
rect 42229 -5729 42419 -5579
rect 47610 -5732 48012 -5580
rect 49233 -5729 49423 -5579
rect 50077 -5729 50093 -5029
rect 50228 -5729 50242 -5029
rect 50077 -8312 50242 -5729
rect 4015 -8636 4215 -8436
rect 11219 -8635 11419 -8435
rect 18423 -8635 18623 -8435
rect 30031 -8634 30231 -8434
rect 37235 -8635 37435 -8435
rect 44439 -8635 44639 -8435
rect 50077 -8651 50082 -8312
rect 50236 -8651 50242 -8312
rect 50077 -8660 50242 -8651
<< via2 >>
rect 50087 26565 50233 26893
rect 50082 -8651 50236 -8312
<< metal3 >>
rect 23355 26554 27812 26904
rect 49400 26893 50261 26904
rect 49400 26565 50087 26893
rect 50233 26565 50261 26893
rect 49400 26554 50261 26565
rect 22121 25941 29057 26341
rect 49400 25941 51288 26341
rect 22121 25341 29057 25741
rect 49400 25341 50667 25741
rect 320 24741 1773 25141
rect 22121 24741 29057 25141
rect 49400 24741 50021 25141
rect 320 -6494 720 24741
rect 889 24141 1773 24541
rect 22121 24141 29057 24541
rect 49400 24141 50021 24541
rect 889 -5894 1289 24141
rect 6971 23990 7774 23992
rect 1451 23810 50052 23990
rect 36772 23690 37012 23691
rect 1451 23510 49752 23690
rect 25478 23360 25629 23510
rect 5891 23160 6091 23360
rect 12895 23160 13095 23360
rect 19899 23160 20099 23360
rect 23554 23164 27683 23360
rect 33907 23160 34107 23360
rect 40911 23160 41111 23360
rect 47915 23160 48115 23360
rect 49572 8332 49752 23510
rect 49872 8827 50052 23810
rect 49871 8731 50052 8827
rect 49852 8531 50052 8731
rect 49552 8132 49753 8332
rect 5891 -5113 6091 -4913
rect 12895 -5113 13095 -4913
rect 19899 -5113 20099 -4913
rect 33907 -5113 34107 -4913
rect 40911 -5113 41111 -4913
rect 47915 -5113 48115 -4913
rect 49572 -5265 49752 8132
rect 1451 -5445 49752 -5265
rect 49872 -5565 50052 8531
rect 1451 -5745 50052 -5565
rect 889 -6294 1775 -5894
rect 22123 -6294 29049 -5894
rect 49402 -6294 50136 -5894
rect 320 -6894 1775 -6494
rect 22123 -6894 29049 -6494
rect 49402 -6894 50136 -6494
rect 50267 -7094 50667 25341
rect 22142 -7494 29058 -7094
rect 49402 -7494 50667 -7094
rect 50888 -7694 51288 25941
rect 22142 -8094 29058 -7694
rect 49402 -8094 51288 -7694
rect 23389 -8657 27796 -8307
rect 49401 -8312 50259 -8306
rect 49401 -8651 50082 -8312
rect 50236 -8651 50259 -8312
rect 49401 -8657 50259 -8651
use EF_AMUX21x  EF_AMUX21x_0
timestamp 1747671550
transform 0 -1 14638 1 0 -9704
box 979 -8763 5769 -1541
use EF_AMUX21x  EF_AMUX21x_1
timestamp 1747671550
transform 0 -1 7434 1 0 -9704
box 979 -8763 5769 -1541
use EF_AMUX21x  x1
timestamp 1747671550
transform 0 -1 26246 -1 0 27951
box 979 -8763 5769 -1541
use EF_AMUX21x  x2
timestamp 1747671550
transform 0 -1 40654 1 0 -9704
box 979 -8763 5769 -1541
use EF_AMUX21x  x3
timestamp 1747671550
transform 0 -1 14638 -1 0 27951
box 979 -8763 5769 -1541
use EF_AMUX21x  x4
timestamp 1747671550
transform 0 -1 7434 -1 0 27951
box 979 -8763 5769 -1541
use EF_AMUX21x  x5
timestamp 1747671550
transform 0 -1 33450 1 0 -9704
box 979 -8763 5769 -1541
use EF_AMUX21x  x8
timestamp 1747671550
transform 0 -1 26246 1 0 -9704
box 979 -8763 5769 -1541
use EF_AMUX21x  x9
timestamp 1747671550
transform 0 -1 230 1 0 -9704
box 979 -8763 5769 -1541
use EF_AMUX21x  x10
timestamp 1747671550
transform 0 -1 40654 -1 0 27951
box 979 -8763 5769 -1541
use EF_AMUX21x  x11
timestamp 1747671550
transform 0 -1 33450 -1 0 27951
box 979 -8763 5769 -1541
use EF_AMUX21x  x12
timestamp 1747671550
transform 0 -1 230 -1 0 27951
box 979 -8763 5769 -1541
<< labels >>
flabel metal3 49852 8531 50052 8731 0 FreeSans 256 180 0 0 VH
port 24 nsew
flabel metal3 49552 8132 49752 8332 0 FreeSans 256 180 0 0 VL
port 25 nsew
flabel metal3 47915 23160 48115 23360 0 FreeSans 256 90 0 0 D5
port 13 nsew
flabel metal3 40911 23160 41111 23360 0 FreeSans 256 90 0 0 D1
port 8 nsew
flabel metal3 33907 23160 34107 23360 0 FreeSans 256 90 0 0 D3
port 2 nsew
flabel metal3 19899 23160 20099 23360 0 FreeSans 256 90 0 0 D8
port 17 nsew
flabel metal3 12895 23160 13095 23360 0 FreeSans 256 90 0 0 D6
port 19 nsew
flabel metal3 5891 23160 6091 23360 0 FreeSans 256 90 0 0 D10
port 27 nsew
flabel metal3 49933 -6220 50133 -6020 0 FreeSans 256 180 0 0 DVSS
port 22 nsew
flabel metal3 49937 -7978 50137 -7778 0 FreeSans 256 180 0 0 VDD
port 20 nsew
flabel metal3 49937 -7385 50137 -7185 0 FreeSans 256 180 0 0 VSS
port 26 nsew
flabel metal3 49935 -6791 50135 -6591 0 FreeSans 256 180 0 0 DVDD
port 21 nsew
flabel metal3 47915 -5113 48115 -4913 0 FreeSans 256 90 0 0 D4
port 10 nsew
flabel metal3 40911 -5113 41111 -4913 0 FreeSans 256 90 0 0 D0
port 5 nsew
flabel metal3 33907 -5113 34107 -4913 0 FreeSans 256 90 0 0 D2
port 0 nsew
flabel metal3 19899 -5113 20099 -4913 0 FreeSans 256 90 0 0 D9
port 15 nsew
flabel metal3 12895 -5113 13095 -4913 0 FreeSans 256 90 0 0 D7
port 18 nsew
flabel metal3 5891 -5113 6091 -4913 0 FreeSans 256 90 0 0 D11
port 28 nsew
flabel metal2 4015 26681 4215 26881 0 FreeSans 256 90 0 0 SELD10
port 29 nsew
flabel metal2 11219 26683 11419 26883 0 FreeSans 256 90 0 0 SELD6
port 16 nsew
flabel metal2 18424 26682 18624 26882 0 FreeSans 256 90 0 0 SELD8
port 12 nsew
flabel metal2 30033 26682 30233 26882 0 FreeSans 256 90 0 0 SELD3
port 3 nsew
flabel metal2 37235 26681 37435 26881 0 FreeSans 256 90 0 0 SELD1
port 6 nsew
flabel metal2 44440 26680 44640 26880 0 FreeSans 256 90 0 0 SELD5
port 9 nsew
flabel metal2 44439 -8635 44639 -8435 0 FreeSans 256 90 0 0 SELD4
port 7 nsew
flabel metal2 37235 -8635 37435 -8435 0 FreeSans 256 90 0 0 SELD0
port 4 nsew
flabel metal2 30031 -8634 30231 -8434 0 FreeSans 256 90 0 0 SELD2
port 1 nsew
flabel metal2 18423 -8635 18623 -8435 0 FreeSans 256 90 0 0 SELD9
port 11 nsew
flabel metal2 11219 -8635 11419 -8435 0 FreeSans 256 90 0 0 SELD7
port 14 nsew
flabel metal2 4015 -8636 4215 -8436 0 FreeSans 256 90 0 0 SELD11
port 30 nsew
flabel metal3 49827 -8586 50026 -8387 0 FreeSans 320 0 0 0 VCM
port 31 nsew
<< properties >>
string MASKHINTS_HVI 49417 -8725 49493 -5254 1705 -8724 1778 -5253 1705 23500 1778 26971 49417 23501 49493 26972
<< end >>
