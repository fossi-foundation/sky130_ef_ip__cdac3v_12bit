magic
tech sky130A
magscale 1 2
timestamp 1747669346
<< error_p >>
rect 66120 -2268 66440 -2244
rect 66120 -2540 66144 -2268
rect 66120 -2564 66440 -2540
rect 66070 -3090 66390 -3066
rect 66070 -3362 66094 -3090
rect 66070 -3386 66390 -3362
<< metal3 >>
rect 66223 -2310 66287 -2304
rect 65895 -2440 66223 -2380
rect 66287 -2434 66288 -2374
rect 66223 -2502 66287 -2496
rect 66223 -3131 66287 -3125
rect 66287 -3251 66615 -3191
rect 66223 -3323 66287 -3317
<< via3 >>
rect 66223 -2496 66287 -2310
rect 66223 -3317 66287 -3131
<< metal4 >>
rect 66225 -2785 66285 -2540
rect 66070 -2845 66440 -2785
rect 66225 -3090 66285 -2845
<< via4 >>
rect 66144 -2310 66416 -2268
rect 66144 -2496 66223 -2310
rect 66223 -2496 66287 -2310
rect 66287 -2496 66416 -2310
rect 66144 -2540 66416 -2496
rect 66094 -3131 66366 -3090
rect 66094 -3317 66223 -3131
rect 66223 -3317 66287 -3131
rect 66287 -3317 66366 -3131
rect 66094 -3362 66366 -3317
<< metal5 >>
rect 66120 -2268 66440 -2244
rect 66120 -2540 66144 -2268
rect 66416 -2540 66440 -2268
rect 66120 -2564 66440 -2540
rect 66070 -3090 66390 -3066
rect 66070 -3362 66094 -3090
rect 66366 -3362 66390 -3090
rect 66070 -3386 66390 -3362
<< end >>
